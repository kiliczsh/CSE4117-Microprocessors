module instreg(inst,clk,A,B,ALU_Sel);
  input inst,clk;
  
  
  
  
  
 endmodule
