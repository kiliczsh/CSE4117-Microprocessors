module instreg(inst,clk,A,B,ALU_Sel);
  input inst,clk;
    output[7:0] A,B;
  output[2:0] ALU_Sel;
  
  
  
  
  
 endmodule
