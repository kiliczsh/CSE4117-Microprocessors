module instreg(inst,clk);
  input inst,clk;
  
  
  
  
 endmodule
