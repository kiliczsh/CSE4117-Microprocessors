module instreg(inst,clk,A,B,ALU_Sel);
  input[7:0] inst;
  input clk;
    output[7:0] A,B;
  output[2:0] ALU_Sel;
  
  
  
  
  
 endmodule
