module datapath();

endmodule
